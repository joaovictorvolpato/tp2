LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY projetofinal IS
PORT (a: IN STD_LOGIC);
END projetofinal;

ARCHITECTURE estrutura OF projetofinal IS
BEGIN
END estrutura;
